module priority_encoder(dout, din, segments,anodes);
output [2:0] dout;
input [7:0] din ;
output [7:0]segments;
output reg [3:0] anodes = 4'b1110;

assign dout = (din[7] ==1'b1 ) ? 3'b111:
(din[6] ==1'b1 ) ? 3'b110:
(din[5] ==1'b1 ) ? 3'b101:
(din[4] ==1'b1) ? 3'b100:
(din[3] ==1'b1) ? 3'b011:
(din[2] ==1'b1) ? 3'b010:
(din[1] ==1'b1) ? 3'b001:
(din[0] ==1'b1) ? 3'b000: 3'bxxx;

segment_decoder uut(.digit(dout),.segments(segments));
endmodule
