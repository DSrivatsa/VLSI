module mult_2_bit(input [1:0]A, input [1:0] B, output reg [3:0] p,output a,b,c,d,e,f,g);
always@(*) begin
p=A*B;
end
assign a=~((p[3])|((p[1])&(p[0]))|((p[2])&(p[0]))|((~(p[2]))&(~(p[0]))));
assign b=~((~(p[2]))|((~(p[1]))&(~(p[0])))|((p[1])&(p[0])));
assign c=~((p[2])|(~(p[1]))|(p[0]));
assign d=~((~(p[2]))&(~(p[0]))|((p[1])&(~(p[0])))|((p[2])&(~(p[1]))&(p[0]))|((~(p[2]))&(p[1])));
assign e=~(((~(p[2]))&(~(p[0])))|((p[1])&(~(p[0]))));
assign f=~((p[3])|((~(p[1]))&(~(p[0])))|((p[2])&(~(p[1])))|((p[2])&(~(p[0]))));
assign g=~((p[3])|((p[2])&(~(p[1])))|((~(p[2]))&(p[1]))|((p[1])&(~(p[0]))));

endmodule
